`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/07/26 19:47:34
// Design Name: 
// Module Name: InstructionMemory
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

//ROM read only memory
//组合逻辑

module InstructionMemory(
    input      [32 -1:0] Address, 
	output reg [32 -1:0] Instruction
    );
always@(*)
begin
//case(Address)
case (Address[10:2])
      9'd0: Instruction<=32'h24080000;	
9'd1: Instruction<=32'h8d100000;	
9'd2: Instruction<=32'h00102021;	
9'd3: Instruction<=32'h21050004;	
9'd4: Instruction<=32'h0c100010;	
9'd5: Instruction<=32'h24080004;	
9'd6: Instruction<=32'h24040000;	
9'd7: Instruction<=32'h3c010010;	
9'd8: Instruction<=32'h34290400;	
9'd9: Instruction<=32'h21290004;	
9'd10: Instruction<=32'h8d2a0000;	
9'd11: Instruction<=32'h008a2020;	
9'd12: Instruction<=32'h21080004;	
9'd13: Instruction<=32'h0106082a;	
9'd14: Instruction<=32'h1420fffa;	
9'd15: Instruction<=32'h0c10003d;	
9'd16: Instruction<=32'h3c010010;	
9'd17: Instruction<=32'h34310400;	
9'd18: Instruction<=32'hae200000;	
9'd19: Instruction<=32'h00043080;	
9'd20: Instruction<=32'h20090001;	
9'd21: Instruction<=32'h200bffff;	
9'd22: Instruction<=32'h00115020;	
9'd23: Instruction<=32'h11240004;	
9'd24: Instruction<=32'h214a0004;	
9'd25: Instruction<=32'had4b0000;	
9'd26: Instruction<=32'h21290001;	
9'd27: Instruction<=32'h1524fffc;	
9'd28: Instruction<=32'h20080001;	
9'd29: Instruction<=32'h00004820;	
9'd30: Instruction<=32'h00005020;	
9'd31: Instruction<=32'h00095940;	
9'd32: Instruction<=32'h016a5820;	
9'd33: Instruction<=32'h02296020;	
9'd34: Instruction<=32'h8d8c0000;	
9'd35: Instruction<=32'h200dffff;	
9'd36: Instruction<=32'h118d000e;	
9'd37: Instruction<=32'h00ab6020;	
9'd38: Instruction<=32'h8d8c0000;	
9'd39: Instruction<=32'h118d000b;	
9'd40: Instruction<=32'h022a7020;	
9'd41: Instruction<=32'h8dce0000;	
9'd42: Instruction<=32'h02297820;	
9'd43: Instruction<=32'h8def0000;	
9'd44: Instruction<=32'h01ec7820;	
9'd45: Instruction<=32'h11cd0003;	
9'd46: Instruction<=32'h01ee082a;	
9'd47: Instruction<=32'h14200001;	
9'd48: Instruction<=32'h08100033;	
9'd49: Instruction<=32'h022a7020;	
9'd50: Instruction<=32'hadcf0000;	
9'd51: Instruction<=32'h214a0004;	
9'd52: Instruction<=32'h0146082a;	
9'd53: Instruction<=32'h1420ffe9;	
9'd54: Instruction<=32'h21290004;	
9'd55: Instruction<=32'h0126082a;	
9'd56: Instruction<=32'h1420ffe5;	
9'd57: Instruction<=32'h21080004;	
9'd58: Instruction<=32'h0106082a;	
9'd59: Instruction<=32'h1420ffe1;	
9'd60: Instruction<=32'h03e00008;	
9'd61: Instruction<=32'h240503e8;	
9'd62: Instruction<=32'h24060000;	
9'd63: Instruction<=32'h3c014000;	
9'd64: Instruction<=32'h34270010;	
9'd65: Instruction<=32'h00044902;	
9'd66: Instruction<=32'h00045202;	
9'd67: Instruction<=32'h00045b02;	
9'd68: Instruction<=32'h3088000f;	
9'd69: Instruction<=32'h3129000f;	
9'd70: Instruction<=32'h314a000f;	
9'd71: Instruction<=32'h316b000f;	
9'd72: Instruction<=32'h15000002;	
9'd73: Instruction<=32'h240c0ec0;	
9'd74: Instruction<=32'hacec0000;	
9'd75: Instruction<=32'h20010001;	
9'd76: Instruction<=32'h14280002;	
9'd77: Instruction<=32'h240c0ef9;	
9'd78: Instruction<=32'hacec0000;	
9'd79: Instruction<=32'h20010002;	
9'd80: Instruction<=32'h14280002;	
9'd81: Instruction<=32'h240c0ea4;	
9'd82: Instruction<=32'hacec0000;	
9'd83: Instruction<=32'h20010003;	
9'd84: Instruction<=32'h14280002;	
9'd85: Instruction<=32'h240c0eb0;	
9'd86: Instruction<=32'hacec0000;	
9'd87: Instruction<=32'h20010004;	
9'd88: Instruction<=32'h14280002;	
9'd89: Instruction<=32'h240c0e99;	
9'd90: Instruction<=32'hacec0000;	
9'd91: Instruction<=32'h20010005;	
9'd92: Instruction<=32'h14280002;	
9'd93: Instruction<=32'h240c0e92;	
9'd94: Instruction<=32'hacec0000;	
9'd95: Instruction<=32'h20010006;	
9'd96: Instruction<=32'h14280002;	
9'd97: Instruction<=32'h240c0e82;	
9'd98: Instruction<=32'hacec0000;	
9'd99: Instruction<=32'h20010007;	
9'd100: Instruction<=32'h14280002;	
9'd101: Instruction<=32'h240c0ef8;	
9'd102: Instruction<=32'hacec0000;	
9'd103: Instruction<=32'h20010008;	
9'd104: Instruction<=32'h14280002;	
9'd105: Instruction<=32'h240c0e80;	
9'd106: Instruction<=32'hacec0000;	
9'd107: Instruction<=32'h20010009;	
9'd108: Instruction<=32'h14280002;	
9'd109: Instruction<=32'h240c0e90;	
9'd110: Instruction<=32'hacec0000;	
9'd111: Instruction<=32'h2001000a;	
9'd112: Instruction<=32'h14280002;	
9'd113: Instruction<=32'h240c0ec8;	
9'd114: Instruction<=32'hacec0000;	
9'd115: Instruction<=32'h2001000b;	
9'd116: Instruction<=32'h14280002;	
9'd117: Instruction<=32'h240c0e83;	
9'd118: Instruction<=32'hacec0000;	
9'd119: Instruction<=32'h2001000c;	
9'd120: Instruction<=32'h14280002;	
9'd121: Instruction<=32'h240c0ec6;	
9'd122: Instruction<=32'hacec0000;	
9'd123: Instruction<=32'h2001000d;	
9'd124: Instruction<=32'h14280002;	
9'd125: Instruction<=32'h240c0ea1;	
9'd126: Instruction<=32'hacec0000;	
9'd127: Instruction<=32'h2001000e;	
9'd128: Instruction<=32'h14280002;	
9'd129: Instruction<=32'h240c0e86;	
9'd130: Instruction<=32'hacec0000;	
9'd131: Instruction<=32'h2001000f;	
9'd132: Instruction<=32'h14280002;	
9'd133: Instruction<=32'h240c0e8e;	
9'd134: Instruction<=32'hacec0000;	
9'd135: Instruction<=32'h20c60001;	
9'd136: Instruction<=32'h14a6ffbf;	
9'd137: Instruction<=32'h00003020;	
9'd138: Instruction<=32'h15200002;	
9'd139: Instruction<=32'h240c0dc0;	
9'd140: Instruction<=32'hacec0000;	
9'd141: Instruction<=32'h20010001;	
9'd142: Instruction<=32'h14290002;	
9'd143: Instruction<=32'h240c0df9;	
9'd144: Instruction<=32'hacec0000;	
9'd145: Instruction<=32'h20010002;	
9'd146: Instruction<=32'h14290002;	
9'd147: Instruction<=32'h240c0da4;	
9'd148: Instruction<=32'hacec0000;	
9'd149: Instruction<=32'h20010003;	
9'd150: Instruction<=32'h14290002;	
9'd151: Instruction<=32'h240c0db0;	
9'd152: Instruction<=32'hacec0000;	
9'd153: Instruction<=32'h20010004;	
9'd154: Instruction<=32'h14290002;	
9'd155: Instruction<=32'h240c0d99;	
9'd156: Instruction<=32'hacec0000;	
9'd157: Instruction<=32'h20010005;	
9'd158: Instruction<=32'h14290002;	
9'd159: Instruction<=32'h240c0d92;	
9'd160: Instruction<=32'hacec0000;	
9'd161: Instruction<=32'h20010006;	
9'd162: Instruction<=32'h14290002;	
9'd163: Instruction<=32'h240c0d82;	
9'd164: Instruction<=32'hacec0000;	
9'd165: Instruction<=32'h20010007;	
9'd166: Instruction<=32'h14290002;	
9'd167: Instruction<=32'h240c0df8;	
9'd168: Instruction<=32'hacec0000;	
9'd169: Instruction<=32'h20010008;	
9'd170: Instruction<=32'h14290002;	
9'd171: Instruction<=32'h240c0d80;	
9'd172: Instruction<=32'hacec0000;	
9'd173: Instruction<=32'h20010009;	
9'd174: Instruction<=32'h14290002;	
9'd175: Instruction<=32'h240c0d90;	
9'd176: Instruction<=32'hacec0000;	
9'd177: Instruction<=32'h2001000a;	
9'd178: Instruction<=32'h14290002;	
9'd179: Instruction<=32'h240c0dc8;	
9'd180: Instruction<=32'hacec0000;	
9'd181: Instruction<=32'h2001000b;	
9'd182: Instruction<=32'h14290002;	
9'd183: Instruction<=32'h240c0d83;	
9'd184: Instruction<=32'hacec0000;	
9'd185: Instruction<=32'h2001000c;	
9'd186: Instruction<=32'h14290002;	
9'd187: Instruction<=32'h240c0dc6;	
9'd188: Instruction<=32'hacec0000;	
9'd189: Instruction<=32'h2001000d;	
9'd190: Instruction<=32'h14290002;	
9'd191: Instruction<=32'h240c0da1;	
9'd192: Instruction<=32'hacec0000;	
9'd193: Instruction<=32'h2001000e;	
9'd194: Instruction<=32'h14290002;	
9'd195: Instruction<=32'h240c0d86;	
9'd196: Instruction<=32'hacec0000;	
9'd197: Instruction<=32'h2001000f;	
9'd198: Instruction<=32'h14290002;	
9'd199: Instruction<=32'h240c0d8e;	
9'd200: Instruction<=32'hacec0000;	
9'd201: Instruction<=32'h20c60001;	
9'd202: Instruction<=32'h14a6ffbf;	
9'd203: Instruction<=32'h00003020;	
9'd204: Instruction<=32'h15400002;	
9'd205: Instruction<=32'h240c0bc0;	
9'd206: Instruction<=32'hacec0000;	
9'd207: Instruction<=32'h20010001;	
9'd208: Instruction<=32'h142a0002;	
9'd209: Instruction<=32'h240c0bf9;	
9'd210: Instruction<=32'hacec0000;	
9'd211: Instruction<=32'h20010002;	
9'd212: Instruction<=32'h142a0002;	
9'd213: Instruction<=32'h240c0ba4;	
9'd214: Instruction<=32'hacec0000;	
9'd215: Instruction<=32'h20010003;	
9'd216: Instruction<=32'h142a0002;	
9'd217: Instruction<=32'h240c0bb0;	
9'd218: Instruction<=32'hacec0000;	
9'd219: Instruction<=32'h20010004;	
9'd220: Instruction<=32'h142a0002;	
9'd221: Instruction<=32'h240c0b99;	
9'd222: Instruction<=32'hacec0000;	
9'd223: Instruction<=32'h20010005;	
9'd224: Instruction<=32'h142a0002;	
9'd225: Instruction<=32'h240c0b92;	
9'd226: Instruction<=32'hacec0000;	
9'd227: Instruction<=32'h20010006;	
9'd228: Instruction<=32'h142a0002;	
9'd229: Instruction<=32'h240c0b82;	
9'd230: Instruction<=32'hacec0000;	
9'd231: Instruction<=32'h20010007;	
9'd232: Instruction<=32'h142a0002;	
9'd233: Instruction<=32'h240c0bf8;	
9'd234: Instruction<=32'hacec0000;	
9'd235: Instruction<=32'h20010008;	
9'd236: Instruction<=32'h142a0002;	
9'd237: Instruction<=32'h240c0b80;	
9'd238: Instruction<=32'hacec0000;	
9'd239: Instruction<=32'h20010009;	
9'd240: Instruction<=32'h142a0002;	
9'd241: Instruction<=32'h240c0b90;	
9'd242: Instruction<=32'hacec0000;	
9'd243: Instruction<=32'h2001000a;	
9'd244: Instruction<=32'h142a0002;	
9'd245: Instruction<=32'h240c0bc8;	
9'd246: Instruction<=32'hacec0000;	
9'd247: Instruction<=32'h2001000b;	
9'd248: Instruction<=32'h142a0002;	
9'd249: Instruction<=32'h240c0b83;	
9'd250: Instruction<=32'hacec0000;	
9'd251: Instruction<=32'h2001000c;	
9'd252: Instruction<=32'h142a0002;	
9'd253: Instruction<=32'h240c0bc6;	
9'd254: Instruction<=32'hacec0000;	
9'd255: Instruction<=32'h2001000d;	
9'd256: Instruction<=32'h142a0002;	
9'd257: Instruction<=32'h240c0ba1;	
9'd258: Instruction<=32'hacec0000;	
9'd259: Instruction<=32'h2001000e;	
9'd260: Instruction<=32'h142a0002;	
9'd261: Instruction<=32'h240c0b86;	
9'd262: Instruction<=32'hacec0000;	
9'd263: Instruction<=32'h2001000f;	
9'd264: Instruction<=32'h142a0002;	
9'd265: Instruction<=32'h240c0b8e;	
9'd266: Instruction<=32'hacec0000;	
9'd267: Instruction<=32'h20c60001;	
9'd268: Instruction<=32'h14a6ffbf;	
9'd269: Instruction<=32'h00003020;	
9'd270: Instruction<=32'h15600002;	
9'd271: Instruction<=32'h240c07c0;	
9'd272: Instruction<=32'hacec0000;	
9'd273: Instruction<=32'h20010001;	
9'd274: Instruction<=32'h142b0002;	
9'd275: Instruction<=32'h240c07f9;	
9'd276: Instruction<=32'hacec0000;	
9'd277: Instruction<=32'h20010002;	
9'd278: Instruction<=32'h142b0002;	
9'd279: Instruction<=32'h240c07a4;	
9'd280: Instruction<=32'hacec0000;	
9'd281: Instruction<=32'h20010003;	
9'd282: Instruction<=32'h142b0002;	
9'd283: Instruction<=32'h240c07b0;	
9'd284: Instruction<=32'hacec0000;	
9'd285: Instruction<=32'h20010004;	
9'd286: Instruction<=32'h142b0002;	
9'd287: Instruction<=32'h240c0799;	
9'd288: Instruction<=32'hacec0000;	
9'd289: Instruction<=32'h20010005;	
9'd290: Instruction<=32'h142b0002;	
9'd291: Instruction<=32'h240c0792;	
9'd292: Instruction<=32'hacec0000;	
9'd293: Instruction<=32'h20010006;	
9'd294: Instruction<=32'h142b0002;	
9'd295: Instruction<=32'h240c0782;	
9'd296: Instruction<=32'hacec0000;	
9'd297: Instruction<=32'h20010007;	
9'd298: Instruction<=32'h142b0002;	
9'd299: Instruction<=32'h240c07f8;	
9'd300: Instruction<=32'hacec0000;	
9'd301: Instruction<=32'h20010008;	
9'd302: Instruction<=32'h142b0002;	
9'd303: Instruction<=32'h240c0780;	
9'd304: Instruction<=32'hacec0000;	
9'd305: Instruction<=32'h20010009;	
9'd306: Instruction<=32'h142b0002;	
9'd307: Instruction<=32'h240c0790;	
9'd308: Instruction<=32'hacec0000;	
9'd309: Instruction<=32'h2001000a;	
9'd310: Instruction<=32'h142b0002;	
9'd311: Instruction<=32'h240c07c8;	
9'd312: Instruction<=32'hacec0000;	
9'd313: Instruction<=32'h2001000b;	
9'd314: Instruction<=32'h142b0002;	
9'd315: Instruction<=32'h240c0783;	
9'd316: Instruction<=32'hacec0000;	
9'd317: Instruction<=32'h2001000c;	
9'd318: Instruction<=32'h142b0002;	
9'd319: Instruction<=32'h240c07c6;	
9'd320: Instruction<=32'hacec0000;	
9'd321: Instruction<=32'h2001000d;	
9'd322: Instruction<=32'h142b0002;	
9'd323: Instruction<=32'h240c07a1;	
9'd324: Instruction<=32'hacec0000;	
9'd325: Instruction<=32'h2001000e;	
9'd326: Instruction<=32'h142b0002;	
9'd327: Instruction<=32'h240c0786;	
9'd328: Instruction<=32'hacec0000;	
9'd329: Instruction<=32'h2001000f;	
9'd330: Instruction<=32'h142b0002;	
9'd331: Instruction<=32'h240c078e;	
9'd332: Instruction<=32'hacec0000;	
9'd333: Instruction<=32'h20c60001;	
9'd334: Instruction<=32'h14a6ffbf;	
9'd335: Instruction<=32'h0810003d;	


        default:Instruction <= 32'h00000000;
endcase
end

endmodule
